module design1(dut_if i);


endmodule
	
	
