
package my_package;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "seq_item.svh"
	`include "sequence.svh"
	`include "driver.svh"
	`include "monitor.svh"
	`include "agent.svh"
	`include "sb.svh"
	`include "environment.svh"
	`include "test.svh"
endpackage
