class base;
	protected int i;
endclass

class ext extends base;
function new();
i=10;
endfunction
endclass
