`timescale 1ns/1ns
package test_pkg ;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "env.svh"
	`include "test.svh"
endpackage 




