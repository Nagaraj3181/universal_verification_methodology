interface dut_if;
 bit clk,rst;
 logic [3:0] count;
endinterface
