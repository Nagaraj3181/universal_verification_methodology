package pack;
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "alu_seq_item.sv"
`include "alu_sequence.sv"
`include "driver.sv"
`include "alu_agent.sv"
`include "env.sv"
`include "test.sv"
endpackage
