package my_pack;
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "transaction.svh"
`include "compa.svh"
`include "cmpb.svh"
`include "env.svh"
`include "test.svh"


endpackage